module axi_2to2_biu (
);




endmodule
