module sram128x64 (
    input               CK,
    input               CS,
    input               WE,
    input        [ 6:0] A,
    input        [ 7:0] BYTE,
    input        [63:0] DI,
    output logic [63:0] DO
);

`ifdef DC
SRAM i_SRAM_0 (
    .A0   ( A[0]         ),
    .A1   ( A[1]         ),
    .A2   ( A[2]         ),
    .A3   ( A[3]         ),
    .A4   ( A[4]         ),
    .A5   ( A[5]         ),
    .A6   ( 1'b0         ),
    .A7   ( 1'b0         ),
    .A8   ( 1'b0         ),
    .A9   ( 1'b0         ),
    .A10  ( 1'b0         ),
    .A11  ( 1'b0         ),
    .A12  ( 1'b0         ),
    .A13  ( 1'b0         ),
    .DO0  ( DO[0]        ),
    .DO1  ( DO[1]        ),
    .DO2  ( DO[2]        ),
    .DO3  ( DO[3]        ),
    .DO4  ( DO[4]        ),
    .DO5  ( DO[5]        ),
    .DO6  ( DO[6]        ),
    .DO7  ( DO[7]        ),
    .DO8  ( DO[8]        ),
    .DO9  ( DO[9]        ),
    .DO10 ( DO[10]       ),
    .DO11 ( DO[11]       ),
    .DO12 ( DO[12]       ),
    .DO13 ( DO[13]       ),
    .DO14 ( DO[14]       ),
    .DO15 ( DO[15]       ),
    .DO16 ( DO[16]       ),
    .DO17 ( DO[17]       ),
    .DO18 ( DO[18]       ),
    .DO19 ( DO[19]       ),
    .DO20 ( DO[20]       ),
    .DO21 ( DO[21]       ),
    .DO22 ( DO[22]       ),
    .DO23 ( DO[23]       ),
    .DO24 ( DO[24]       ),
    .DO25 ( DO[25]       ),
    .DO26 ( DO[26]       ),
    .DO27 ( DO[27]       ),
    .DO28 ( DO[28]       ),
    .DO29 ( DO[29]       ),
    .DO30 ( DO[30]       ),
    .DO31 ( DO[31]       ),
    .DI0  ( DI[0]        ),
    .DI1  ( DI[1]        ),
    .DI2  ( DI[2]        ),
    .DI3  ( DI[3]        ),
    .DI4  ( DI[4]        ),
    .DI5  ( DI[5]        ),
    .DI6  ( DI[6]        ),
    .DI7  ( DI[7]        ),
    .DI8  ( DI[8]        ),
    .DI9  ( DI[9]        ),
    .DI10 ( DI[10]       ),
    .DI11 ( DI[11]       ),
    .DI12 ( DI[12]       ),
    .DI13 ( DI[13]       ),
    .DI14 ( DI[14]       ),
    .DI15 ( DI[15]       ),
    .DI16 ( DI[16]       ),
    .DI17 ( DI[17]       ),
    .DI18 ( DI[18]       ),
    .DI19 ( DI[19]       ),
    .DI20 ( DI[20]       ),
    .DI21 ( DI[21]       ),
    .DI22 ( DI[22]       ),
    .DI23 ( DI[23]       ),
    .DI24 ( DI[24]       ),
    .DI25 ( DI[25]       ),
    .DI26 ( DI[26]       ),
    .DI27 ( DI[27]       ),
    .DI28 ( DI[28]       ),
    .DI29 ( DI[29]       ),
    .DI30 ( DI[30]       ),
    .DI31 ( DI[31]       ),
    .CK   ( CK           ),
    .WEB0 ( ~BYTE[0]     ),
    .WEB1 ( ~BYTE[1]     ),
    .WEB2 ( ~BYTE[2]     ),
    .WEB3 ( ~BYTE[3]     ),
    .OE   ( 1'b1         ),
    .CS   ( CS           )
);
SRAM i_SRAM_1 (
    .A0   ( A[0]         ),
    .A1   ( A[1]         ),
    .A2   ( A[2]         ),
    .A3   ( A[3]         ),
    .A4   ( A[4]         ),
    .A5   ( A[5]         ),
    .A6   ( 1'b0         ),
    .A7   ( 1'b0         ),
    .A8   ( 1'b0         ),
    .A9   ( 1'b0         ),
    .A10  ( 1'b0         ),
    .A11  ( 1'b0         ),
    .A12  ( 1'b0         ),
    .A13  ( 1'b0         ),
    .DO0  ( DO[32+0]     ),
    .DO1  ( DO[32+1]     ),
    .DO2  ( DO[32+2]     ),
    .DO3  ( DO[32+3]     ),
    .DO4  ( DO[32+4]     ),
    .DO5  ( DO[32+5]     ),
    .DO6  ( DO[32+6]     ),
    .DO7  ( DO[32+7]     ),
    .DO8  ( DO[32+8]     ),
    .DO9  ( DO[32+9]     ),
    .DO10 ( DO[32+10]    ),
    .DO11 ( DO[32+11]    ),
    .DO12 ( DO[32+12]    ),
    .DO13 ( DO[32+13]    ),
    .DO14 ( DO[32+14]    ),
    .DO15 ( DO[32+15]    ),
    .DO16 ( DO[32+16]    ),
    .DO17 ( DO[32+17]    ),
    .DO18 ( DO[32+18]    ),
    .DO19 ( DO[32+19]    ),
    .DO20 ( DO[32+20]    ),
    .DO21 ( DO[32+21]    ),
    .DO22 ( DO[32+22]    ),
    .DO23 ( DO[32+23]    ),
    .DO24 ( DO[32+24]    ),
    .DO25 ( DO[32+25]    ),
    .DO26 ( DO[32+26]    ),
    .DO27 ( DO[32+27]    ),
    .DO28 ( DO[32+28]    ),
    .DO29 ( DO[32+29]    ),
    .DO30 ( DO[32+30]    ),
    .DO31 ( DO[32+31]    ),
    .DI0  ( DI[32+0]     ),
    .DI1  ( DI[32+1]     ),
    .DI2  ( DI[32+2]     ),
    .DI3  ( DI[32+3]     ),
    .DI4  ( DI[32+4]     ),
    .DI5  ( DI[32+5]     ),
    .DI6  ( DI[32+6]     ),
    .DI7  ( DI[32+7]     ),
    .DI8  ( DI[32+8]     ),
    .DI9  ( DI[32+9]     ),
    .DI10 ( DI[32+10]    ),
    .DI11 ( DI[32+11]    ),
    .DI12 ( DI[32+12]    ),
    .DI13 ( DI[32+13]    ),
    .DI14 ( DI[32+14]    ),
    .DI15 ( DI[32+15]    ),
    .DI16 ( DI[32+16]    ),
    .DI17 ( DI[32+17]    ),
    .DI18 ( DI[32+18]    ),
    .DI19 ( DI[32+19]    ),
    .DI20 ( DI[32+20]    ),
    .DI21 ( DI[32+21]    ),
    .DI22 ( DI[32+22]    ),
    .DI23 ( DI[32+23]    ),
    .DI24 ( DI[32+24]    ),
    .DI25 ( DI[32+25]    ),
    .DI26 ( DI[32+26]    ),
    .DI27 ( DI[32+27]    ),
    .DI28 ( DI[32+28]    ),
    .DI29 ( DI[32+29]    ),
    .DI30 ( DI[32+30]    ),
    .DI31 ( DI[32+31]    ),
    .CK   ( CK           ),
    .WEB0 ( ~BYTE[4+0]   ),
    .WEB1 ( ~BYTE[4+1]   ),
    .WEB2 ( ~BYTE[4+2]   ),
    .WEB3 ( ~BYTE[4+3]   ),
    .OE   ( 1'b1         ),
    .CS   ( CS           )
);
SRAM i_SRAM_2 (
    .A0   ( A[0]         ),
    .A1   ( A[1]         ),
    .A2   ( A[2]         ),
    .A3   ( A[3]         ),
    .A4   ( A[4]         ),
    .A5   ( A[5]         ),
    .A6   ( 1'b0         ),
    .A7   ( 1'b0         ),
    .A8   ( 1'b0         ),
    .A9   ( 1'b0         ),
    .A10  ( 1'b0         ),
    .A11  ( 1'b0         ),
    .A12  ( 1'b0         ),
    .A13  ( 1'b0         ),
    .DO0  ( DO[64+0]     ),
    .DO1  ( DO[64+1]     ),
    .DO2  ( DO[64+2]     ),
    .DO3  ( DO[64+3]     ),
    .DO4  ( DO[64+4]     ),
    .DO5  ( DO[64+5]     ),
    .DO6  ( DO[64+6]     ),
    .DO7  ( DO[64+7]     ),
    .DO8  ( DO[64+8]     ),
    .DO9  ( DO[64+9]     ),
    .DO10 ( DO[64+10]    ),
    .DO11 ( DO[64+11]    ),
    .DO12 ( DO[64+12]    ),
    .DO13 ( DO[64+13]    ),
    .DO14 ( DO[64+14]    ),
    .DO15 ( DO[64+15]    ),
    .DO16 ( DO[64+16]    ),
    .DO17 ( DO[64+17]    ),
    .DO18 ( DO[64+18]    ),
    .DO19 ( DO[64+19]    ),
    .DO20 ( DO[64+20]    ),
    .DO21 ( DO[64+21]    ),
    .DO22 ( DO[64+22]    ),
    .DO23 ( DO[64+23]    ),
    .DO24 ( DO[64+24]    ),
    .DO25 ( DO[64+25]    ),
    .DO26 ( DO[64+26]    ),
    .DO27 ( DO[64+27]    ),
    .DO28 ( DO[64+28]    ),
    .DO29 ( DO[64+29]    ),
    .DO30 ( DO[64+30]    ),
    .DO31 ( DO[64+31]    ),
    .DI0  ( DI[64+0]     ),
    .DI1  ( DI[64+1]     ),
    .DI2  ( DI[64+2]     ),
    .DI3  ( DI[64+3]     ),
    .DI4  ( DI[64+4]     ),
    .DI5  ( DI[64+5]     ),
    .DI6  ( DI[64+6]     ),
    .DI7  ( DI[64+7]     ),
    .DI8  ( DI[64+8]     ),
    .DI9  ( DI[64+9]     ),
    .DI10 ( DI[64+10]    ),
    .DI11 ( DI[64+11]    ),
    .DI12 ( DI[64+12]    ),
    .DI13 ( DI[64+13]    ),
    .DI14 ( DI[64+14]    ),
    .DI15 ( DI[64+15]    ),
    .DI16 ( DI[64+16]    ),
    .DI17 ( DI[64+17]    ),
    .DI18 ( DI[64+18]    ),
    .DI19 ( DI[64+19]    ),
    .DI20 ( DI[64+20]    ),
    .DI21 ( DI[64+21]    ),
    .DI22 ( DI[64+22]    ),
    .DI23 ( DI[64+23]    ),
    .DI24 ( DI[64+24]    ),
    .DI25 ( DI[64+25]    ),
    .DI26 ( DI[64+26]    ),
    .DI27 ( DI[64+27]    ),
    .DI28 ( DI[64+28]    ),
    .DI29 ( DI[64+29]    ),
    .DI30 ( DI[64+30]    ),
    .DI31 ( DI[64+31]    ),
    .CK   ( CK           ),
    .WEB0 ( ~BYTE[8+0]   ),
    .WEB1 ( ~BYTE[8+1]   ),
    .WEB2 ( ~BYTE[8+2]   ),
    .WEB3 ( ~BYTE[8+3]   ),
    .OE   ( 1'b1         ),
    .CS   ( CS           )
);
SRAM i_SRAM_3 (
    .A0   ( A[0]         ),
    .A1   ( A[1]         ),
    .A2   ( A[2]         ),
    .A3   ( A[3]         ),
    .A4   ( A[4]         ),
    .A5   ( A[5]         ),
    .A6   ( 1'b0         ),
    .A7   ( 1'b0         ),
    .A8   ( 1'b0         ),
    .A9   ( 1'b0         ),
    .A10  ( 1'b0         ),
    .A11  ( 1'b0         ),
    .A12  ( 1'b0         ),
    .A13  ( 1'b0         ),
    .DO0  ( DO[96+0]     ),
    .DO1  ( DO[96+1]     ),
    .DO2  ( DO[96+2]     ),
    .DO3  ( DO[96+3]     ),
    .DO4  ( DO[96+4]     ),
    .DO5  ( DO[96+5]     ),
    .DO6  ( DO[96+6]     ),
    .DO7  ( DO[96+7]     ),
    .DO8  ( DO[96+8]     ),
    .DO9  ( DO[96+9]     ),
    .DO10 ( DO[96+10]    ),
    .DO11 ( DO[96+11]    ),
    .DO12 ( DO[96+12]    ),
    .DO13 ( DO[96+13]    ),
    .DO14 ( DO[96+14]    ),
    .DO15 ( DO[96+15]    ),
    .DO16 ( DO[96+16]    ),
    .DO17 ( DO[96+17]    ),
    .DO18 ( DO[96+18]    ),
    .DO19 ( DO[96+19]    ),
    .DO20 ( DO[96+20]    ),
    .DO21 ( DO[96+21]    ),
    .DO22 ( DO[96+22]    ),
    .DO23 ( DO[96+23]    ),
    .DO24 ( DO[96+24]    ),
    .DO25 ( DO[96+25]    ),
    .DO26 ( DO[96+26]    ),
    .DO27 ( DO[96+27]    ),
    .DO28 ( DO[96+28]    ),
    .DO29 ( DO[96+29]    ),
    .DO30 ( DO[96+30]    ),
    .DO31 ( DO[96+31]    ),
    .DI0  ( DI[96+0]     ),
    .DI1  ( DI[96+1]     ),
    .DI2  ( DI[96+2]     ),
    .DI3  ( DI[96+3]     ),
    .DI4  ( DI[96+4]     ),
    .DI5  ( DI[96+5]     ),
    .DI6  ( DI[96+6]     ),
    .DI7  ( DI[96+7]     ),
    .DI8  ( DI[96+8]     ),
    .DI9  ( DI[96+9]     ),
    .DI10 ( DI[96+10]    ),
    .DI11 ( DI[96+11]    ),
    .DI12 ( DI[96+12]    ),
    .DI13 ( DI[96+13]    ),
    .DI14 ( DI[96+14]    ),
    .DI15 ( DI[96+15]    ),
    .DI16 ( DI[96+16]    ),
    .DI17 ( DI[96+17]    ),
    .DI18 ( DI[96+18]    ),
    .DI19 ( DI[96+19]    ),
    .DI20 ( DI[96+20]    ),
    .DI21 ( DI[96+21]    ),
    .DI22 ( DI[96+22]    ),
    .DI23 ( DI[96+23]    ),
    .DI24 ( DI[96+24]    ),
    .DI25 ( DI[96+25]    ),
    .DI26 ( DI[96+26]    ),
    .DI27 ( DI[96+27]    ),
    .DI28 ( DI[96+28]    ),
    .DI29 ( DI[96+29]    ),
    .DI30 ( DI[96+30]    ),
    .DI31 ( DI[96+31]    ),
    .CK   ( CK           ),
    .WEB0 ( ~BYTE[12+0]  ),
    .WEB1 ( ~BYTE[12+1]  ),
    .WEB2 ( ~BYTE[12+2]  ),
    .WEB3 ( ~BYTE[12+3]  ),
    .OE   ( 1'b1         ),
    .CS   ( CS           )
);
`else
logic [63:0] data_out_pre;
logic [63:0] memory [128];

assign data_out_pre = CS ? memory[A] : 64'hx;

always_ff @(posedge CK) begin
    integer i;

    if (CS & WE) begin
        for (i = 0; i < 8; i = i + 1) begin
            if (BYTE[i]) memory[A][i*8+:8] <= DI[i*8+:8];
        end
    end
end

always_ff @(posedge CK) begin
    DO <= data_out_pre;
end
`endif

endmodule
