parameter [`CSR_OP_LEN - 1:0] CSR_OP_NONE = `CSR_OP_LEN'b00,
                              CSR_OP_SET  = `CSR_OP_LEN'b01,
                              CSR_OP_CLR  = `CSR_OP_LEN'b10;
