`define JALR(RS1) {12'b0, RS1, 3'b000, 5'b00000, 7'b1100111}
`define ADDI(RD, RS1, IMM) {IMM, RS1, 3'b000, RD, 7'b0010011}

initial begin
    repeat (100) @(negedge clk);
    dbgapb_wr(`DBGAPB_DBG_EN, 32'b1);
    dbgapb_wr(`DBGAPB_INST, {20'b0, `INST_ATTACH});
    dbgapb_wr(`DBGAPB_INST_WR, 32'b1);
    dbg_rdata = `XLEN'b0;
    dbgapb_status_rd;
    while (dbg_rdata != `XLEN'h3) begin
        @(negedge clk);
        dbgapb_status_rd;
    end
    dbgapb_pc_rd;
    dbgapb_exec(`ADDI(`GPR_T0_ADDR, `GPR_ZERO_ADDR, 12'hcc));
    dbgapb_exec(`JALR(`GPR_T0_ADDR));
    dbgapb_pc_rd;
    dbgapb_pc_rd;
    dbgapb_pc_rd;
    dbgapb_gpr_rd(5'h0);
    dbgapb_gpr_rd(5'h1);
    dbgapb_gpr_rd(5'h2);
    dbgapb_gpr_rd(5'h3);
    dbgapb_gpr_rd(5'h4);
    dbgapb_gpr_rd(5'h5);
    dbgapb_gpr_rd(5'h6);
    dbgapb_gpr_rd(5'h7);
    dbgapb_gpr_rd(5'h8);
    dbgapb_gpr_rd(5'h9);
    dbgapb_gpr_rd(5'ha);
    dbgapb_gpr_rd(5'hb);
    dbgapb_gpr_rd(5'hc);
    dbgapb_gpr_rd(5'hd);
    dbgapb_gpr_rd(5'he);
    dbgapb_gpr_rd(5'hf);
    dbgapb_gpr_rd(5'h10);
    dbgapb_gpr_rd(5'h11);
    dbgapb_gpr_rd(5'h12);
    dbgapb_gpr_rd(5'h13);
    dbgapb_gpr_rd(5'h14);
    dbgapb_gpr_rd(5'h15);
    dbgapb_gpr_rd(5'h16);
    dbgapb_gpr_rd(5'h17);
    dbgapb_gpr_rd(5'h18);
    dbgapb_gpr_rd(5'h19);
    dbgapb_gpr_rd(5'h1a);
    dbgapb_gpr_rd(5'h1b);
    dbgapb_gpr_rd(5'h1c);
    dbgapb_gpr_rd(5'h1d);
    dbgapb_gpr_rd(5'h1e);
    dbgapb_gpr_rd(5'h1f);
    dbgapb_gpr_wr(5'h0 , {32'h0 , 32'h0 });
    dbgapb_gpr_wr(5'h1 , {32'h1 , 32'h1 });
    dbgapb_gpr_wr(5'h2 , {32'h2 , 32'h2 });
    dbgapb_gpr_wr(5'h3 , {32'h3 , 32'h3 });
    dbgapb_gpr_wr(5'h4 , {32'h4 , 32'h4 });
    dbgapb_gpr_wr(5'h5 , {32'h5 , 32'h5 });
    dbgapb_gpr_wr(5'h6 , {32'h6 , 32'h6 });
    dbgapb_gpr_wr(5'h7 , {32'h7 , 32'h7 });
    dbgapb_gpr_wr(5'h8 , {32'h8 , 32'h8 });
    dbgapb_gpr_wr(5'h9 , {32'h9 , 32'h9 });
    dbgapb_gpr_wr(5'ha , {32'ha , 32'ha });
    dbgapb_gpr_wr(5'hb , {32'hb , 32'hb });
    dbgapb_gpr_wr(5'hc , {32'hc , 32'hc });
    dbgapb_gpr_wr(5'hd , {32'hd , 32'hd });
    dbgapb_gpr_wr(5'he , {32'he , 32'he });
    dbgapb_gpr_wr(5'hf , {32'hf , 32'hf });
    dbgapb_gpr_wr(5'h10, {32'h10, 32'h10});
    dbgapb_gpr_wr(5'h11, {32'h11, 32'h11});
    dbgapb_gpr_wr(5'h12, {32'h12, 32'h12});
    dbgapb_gpr_wr(5'h13, {32'h13, 32'h13});
    dbgapb_gpr_wr(5'h14, {32'h14, 32'h14});
    dbgapb_gpr_wr(5'h15, {32'h15, 32'h15});
    dbgapb_gpr_wr(5'h16, {32'h16, 32'h16});
    dbgapb_gpr_wr(5'h17, {32'h17, 32'h17});
    dbgapb_gpr_wr(5'h18, {32'h18, 32'h18});
    dbgapb_gpr_wr(5'h19, {32'h19, 32'h19});
    dbgapb_gpr_wr(5'h1a, {32'h1a, 32'h1a});
    dbgapb_gpr_wr(5'h1b, {32'h1b, 32'h1b});
    dbgapb_gpr_wr(5'h1c, {32'h1c, 32'h1c});
    dbgapb_gpr_wr(5'h1d, {32'h1d, 32'h1d});
    dbgapb_gpr_wr(5'h1e, {32'h1e, 32'h1e});
    dbgapb_gpr_wr(5'h1f, {32'h1f, 32'h1f});
    dbgapb_gpr_rd(5'h0);
    dbgapb_gpr_rd(5'h1);
    dbgapb_gpr_rd(5'h2);
    dbgapb_gpr_rd(5'h3);
    dbgapb_gpr_rd(5'h4);
    dbgapb_gpr_rd(5'h5);
    dbgapb_gpr_rd(5'h6);
    dbgapb_gpr_rd(5'h7);
    dbgapb_gpr_rd(5'h8);
    dbgapb_gpr_rd(5'h9);
    dbgapb_gpr_rd(5'ha);
    dbgapb_gpr_rd(5'hb);
    dbgapb_gpr_rd(5'hc);
    dbgapb_gpr_rd(5'hd);
    dbgapb_gpr_rd(5'he);
    dbgapb_gpr_rd(5'hf);
    dbgapb_gpr_rd(5'h10);
    dbgapb_gpr_rd(5'h11);
    dbgapb_gpr_rd(5'h12);
    dbgapb_gpr_rd(5'h13);
    dbgapb_gpr_rd(5'h14);
    dbgapb_gpr_rd(5'h15);
    dbgapb_gpr_rd(5'h16);
    dbgapb_gpr_rd(5'h17);
    dbgapb_gpr_rd(5'h18);
    dbgapb_gpr_rd(5'h19);
    dbgapb_gpr_rd(5'h1a);
    dbgapb_gpr_rd(5'h1b);
    dbgapb_gpr_rd(5'h1c);
    dbgapb_gpr_rd(5'h1d);
    dbgapb_gpr_rd(5'h1e);
    dbgapb_gpr_rd(5'h1f);
    dbgapb_csr_rd(12'h300);
    dbgapb_csr_wr(12'h300, 64'hffffffff_ffffffff);
    dbgapb_csr_rd(12'h300);
    dbgapb_exec(`ADDI(`GPR_ZERO_ADDR, `GPR_ZERO_ADDR, 12'h000));
    dbgapb_wr(`DBGAPB_INST, {20'b0, `INST_RESUME});
    dbgapb_wr(`DBGAPB_INST_WR, 32'b1);
end
