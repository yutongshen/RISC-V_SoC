parameter [2:0] FUNCT3_JALR    = 3'b000,
                FUNCT3_BEQ     = 3'b000,
                FUNCT3_BNE     = 3'b001,
                FUNCT3_BLT     = 3'b100,
                FUNCT3_BGE     = 3'b101,
                FUNCT3_BLTU    = 3'b110,
                FUNCT3_BGEU    = 3'b111,
                FUNCT3_LB      = 3'b000,
                FUNCT3_LH      = 3'b001,
                FUNCT3_LW      = 3'b010,
                FUNCT3_LD      = 3'b011,
                FUNCT3_LBU     = 3'b100,
                FUNCT3_LHU     = 3'b101,
                FUNCT3_LWU     = 3'b110,
                FUNCT3_SB      = 3'b000,
                FUNCT3_SH      = 3'b001,
                FUNCT3_SW      = 3'b010,
                FUNCT3_SD      = 3'b011,
                FUNCT3_ADDI    = 3'b000,
                FUNCT3_SLTI    = 3'b010,
                FUNCT3_SLTIU   = 3'b011,
                FUNCT3_XORI    = 3'b100,
                FUNCT3_ORI     = 3'b110,
                FUNCT3_ANDI    = 3'b111,
                FUNCT3_SLLI    = 3'b001,
                FUNCT3_SRLI    = 3'b101,
                FUNCT3_SRAI    = 3'b101,
                FUNCT3_ADD     = 3'b000,
                FUNCT3_SUB     = 3'b000,
                FUNCT3_SLL     = 3'b001,
                FUNCT3_SLT     = 3'b010,
                FUNCT3_SLTU    = 3'b011,
                FUNCT3_XOR     = 3'b100,
                FUNCT3_SRL     = 3'b101,
                FUNCT3_SRA     = 3'b101,
                FUNCT3_OR      = 3'b110,
                FUNCT3_AND     = 3'b111,
                FUNCT3_FENCE   = 3'b000,
                FUNCT3_FENCE_I = 3'b001,
                FUNCT3_PRIV    = 3'b000,
                FUNCT3_CSRRW   = 3'b001,
                FUNCT3_CSRRS   = 3'b010,
                FUNCT3_CSRRC   = 3'b011,
                FUNCT3_CSRRWI  = 3'b101,
                FUNCT3_CSRRSI  = 3'b110,
                FUNCT3_CSRRCI  = 3'b111,
                FUNCT3_MUL     = 3'b000,
                FUNCT3_MULH    = 3'b001,
                FUNCT3_MULHSU  = 3'b010,
                FUNCT3_MULHU   = 3'b011,
                FUNCT3_DIV     = 3'b100,
                FUNCT3_DIVU    = 3'b101,
                FUNCT3_REM     = 3'b110,
                FUNCT3_REMU    = 3'b111;

parameter [4:0] FUNCT5_LR      = 5'b00010,
                FUNCT5_SC      = 5'b00011,
                FUNCT5_AMOSWAP = 5'b00001,
                FUNCT5_AMOADD  = 5'b00000,
                FUNCT5_AMOXOR  = 5'b00100,
                FUNCT5_AMOAND  = 5'b01100,
                FUNCT5_AMOOR   = 5'b01000,
                FUNCT5_AMOMIN  = 5'b10000,
                FUNCT5_AMOMAX  = 5'b10100,
                FUNCT5_AMOMINU = 5'b11000,
                FUNCT5_AMOMAXU = 5'b11100;

parameter [6:0] FUNCT7_SLLI       = 7'b0000000,
                FUNCT7_SRLI       = 7'b0000000,
                FUNCT7_SRAI       = 7'b0100000,
                FUNCT7_OP0        = 7'b0000000,
                FUNCT7_OP1        = 7'b0100000,
                FUNCT7_SFENCE_VMA = 7'b0001001,
                FUNCT7_MULDIV     = 7'b0000001;

parameter [11:0] FUNCT12_ECALL  = 12'h000,
                 FUNCT12_EBREAK = 12'h001,
                 FUNCT12_WFI    = 12'h105,
                 FUNCT12_SRET   = 12'h102,
                 FUNCT12_MRET   = 12'h302;

// RVC
parameter [2:0] FUNCT3_C0_ADDI4SPN = 3'b000,
                FUNCT3_C0_FLD      = 3'b001,
                FUNCT3_C0_LW       = 3'b010,
                FUNCT3_C0_FLW      = 3'b011,
                FUNCT3_C0_FSD      = 3'b101,
                FUNCT3_C0_SW       = 3'b110,
                FUNCT3_C0_FSW      = 3'b111;

parameter [2:0] FUNCT3_C1_ADDI     = 3'b000,
                FUNCT3_C1_JAL      = 3'b001,
                FUNCT3_C1_LI       = 3'b010,
                FUNCT3_C1_LUI      = 3'b011,
                FUNCT3_C1_OP       = 3'b100,
                FUNCT3_C1_J        = 3'b101,
                FUNCT3_C1_BEQZ     = 3'b110,
                FUNCT3_C1_BNEZ     = 3'b111;

parameter [2:0] FUNCT3_C2_SLLI     = 3'b000,
                FUNCT3_C2_FLDSP    = 3'b001,
                FUNCT3_C2_LWSP     = 3'b010,
                FUNCT3_C2_FLWSP    = 3'b011,
                FUNCT3_C2_OP       = 3'b100,
                FUNCT3_C2_FSDSP    = 3'b101,
                FUNCT3_C2_SWSP     = 3'b110,
                FUNCT3_C2_FSWSP    = 3'b111;

parameter [2:0] FUNCT2_OP_IMM_C_SRLI = 2'b00,
                FUNCT2_OP_IMM_C_SRAI = 2'b01,
                FUNCT2_OP_IMM_C_ANDI = 2'b10,
                FUNCT2_OP_IMM_C_OP   = 2'b11;

parameter [2:0] FUNCT2_OP_C_SUB  = 2'b00,
                FUNCT2_OP_C_XOR  = 2'b01,
                FUNCT2_OP_C_OR   = 2'b10,
                FUNCT2_OP_C_AND  = 2'b11,
                FUNCT2_OP_C_SUBW = 2'b00,
                FUNCT2_OP_C_ADDW = 2'b01;
