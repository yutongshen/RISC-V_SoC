parameter [`BPU_OP_LEN - 1:0] BPU_EQ  = `BPU_OP_LEN'b00,
                              BPU_LT  = `BPU_OP_LEN'b01,
                              BPU_LTU = `BPU_OP_LEN'b10;
